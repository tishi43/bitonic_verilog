//--------------------------------------------------------------------------------------------------
// Copyright (C) 2013-2017 qiu bin 
// All rights reserved   
// Design    : bitstream_p
// Author(s) : qiu bin
// Email     : chat1@126.com
// Phone 15957074161
// QQ:1517642772             
//-------------------------------------------------------------------------------------------------



// used for storing intra4x4_pred_mode, ref_idx, mvp etc
// 
module ram_simple_dual
(
clk,
en,
we,
addra,
addrb,
dia,
dob
);

parameter addr_bits = 7;
parameter data_bits = 100;
input     clk;
input     en;
input     we;
input     [addr_bits-1:0]  addra;
input     [addr_bits-1:0]  addrb;
input     [data_bits-1:0]  dia;
output    [data_bits-1:0]  dob;

wire      clk;
wire      en;
wire      we;
wire      [addr_bits-1:0]  addra;
wire      [addr_bits-1:0]  addrb;
wire      [data_bits-1:0]  dia;
reg       [data_bits-1:0]  dob;

(* ram_style = "block" *)
reg       [data_bits-1:0]  ram[0:(1 << addr_bits) -1];

wire      [data_bits/2-1:0] data[0:(1<<(addr_bits+1))-1];

assign data = ram;

initial  begin
    /*ram = {{50'd38,50'd113},{50'd190,50'd170},{50'd246,50'd177},{50'd111,50'd186},{50'd79,50'd251},{50'd2,50'd121},{50'd91,50'd185},{50'd90,50'd112},
           {50'd132,50'd219},{50'd95,50'd204},{50'd205,50'd69},{50'd54,50'd237},{50'd81,50'd172},{50'd143,50'd138},{50'd18,50'd33},{50'd43,50'd224},
           {50'd244,50'd117},{50'd217,50'd86},{50'd247,50'd24},{50'd83,50'd10},{50'd230,50'd124},{50'd200,50'd233},{50'd151,50'd136},{50'd46,50'd122},
           {50'd85,50'd181},{50'd127,50'd131},{50'd70,50'd14},{50'd254,50'd163},{50'd249,50'd213},{50'd30,50'd193},{50'd13,50'd120},{50'd212,50'd128},
           {50'd32,50'd137},{50'd201,50'd65},{50'd40,50'd116},{50'd159,50'd144},{50'd142,50'd28},{50'd73,50'd240},{50'd236,50'd75},{50'd68,50'd102},
           {50'd4,50'd45},{50'd103,50'd64},{50'd108,50'd179},{50'd243,50'd92},{50'd55,50'd169},{50'd98,50'd182},{50'd82,50'd106},{50'd234,50'd168},
           {50'd44,50'd6},{50'd0,50'd20},{50'd175,50'd80},{50'd135,50'd52},{50'd62,50'd61},{50'd198,50'd199},{50'd166,50'd145},{50'd133,50'd150},
           {50'd51,50'd100},{50'd214,50'd97},{50'd148,50'd192},{50'd149,50'd84},{50'd58,50'd180},{50'd223,50'd250},{50'd130,50'd25},{50'd63,50'd114},
           {50'd160,50'd94},{50'd245,50'd229},{50'd49,50'd16},{50'd50,50'd253},{50'd152,50'd207},{50'd206,50'd5},{50'd203,50'd48},{50'd140,50'd53},
           {50'd57,50'd35},{50'd1,50'd42},{50'd27,50'd71},{50'd156,50'd154},{50'd157,50'd216},{50'd232,50'd239},{50'd218,50'd56},{50'd118,50'd15},
           {50'd29,50'd184},{50'd26,50'd76},{50'd12,50'd99},{50'd155,50'd89},{50'd36,50'd109},{50'd176,50'd255},{50'd72,50'd252},{50'd221,50'd248},
           {50'd197,50'd8},{50'd183,50'd134},{50'd195,50'd226},{50'd66,50'd141},{50'd104,50'd125},{50'd88,50'd209},{50'd194,50'd235},{50'd96,50'd119},
           {50'd202,50'd105},{50'd164,50'd227},{50'd7,50'd208},{50'd123,50'd189},{50'd241,50'd196},{50'd210,50'd74},{50'd3,50'd174},{50'd173,50'd37},
           {50'd21,50'd187},{50'd77,50'd220},{50'd78,50'd87},{50'd191,50'd161},{50'd31,50'd129},{50'd147,50'd19},{50'd93,50'd22},{50'd211,50'd165},
           {50'd23,50'd126},{50'd110,50'd146},{50'd171,50'd167},{50'd242,50'd139},{50'd158,50'd153},{50'd59,50'd34},{50'd67,50'd222},{50'd115,50'd231},
           {50'd39,50'd9},{50'd101,50'd60},{50'd47,50'd215},{50'd178,50'd11},{50'd228,50'd225},{50'd17,50'd162},{50'd238,50'd188},{50'd41,50'd107}};*/


ram = {{50'd252,50'd2040},{50'd700,50'd100},{50'd609,50'd548},{50'd692,50'd1454},{50'd1646,50'd1041},{50'd1923,50'd155},{50'd72,50'd311},{50'd1957,50'd56},
        {50'd1713,50'd1334},{50'd517,50'd381},{50'd1086,50'd980},{50'd1502,50'd14},{50'd375,50'd1944},{50'd550,50'd780},{50'd575,50'd1741},{50'd128,50'd341},
        {50'd1082,50'd1294},{50'd1677,50'd405},{50'd333,50'd561},{50'd1503,50'd1684},{50'd1034,50'd204},{50'd839,50'd479},{50'd1316,50'd1447},{50'd1442,50'd221},
        {50'd1599,50'd1087},{50'd1192,50'd1367},{50'd1196,50'd1515},{50'd1904,50'd642},{50'd940,50'd872},{50'd1623,50'd643},{50'd713,50'd1767},{50'd929,50'd636},
        {50'd345,50'd314},{50'd1702,50'd1962},{50'd1410,50'd429},{50'd1851,50'd419},{50'd459,50'd1012},{50'd1840,50'd555},{50'd1326,50'd815},{50'd1349,50'd151},
        {50'd1016,50'd641},{50'd332,50'd1009},{50'd105,50'd348},{50'd1135,50'd695},{50'd2044,50'd1803},{50'd1364,50'd1968},{50'd1417,50'd264},{50'd958,50'd1037},
        {50'd1894,50'd46},{50'd725,50'd1789},{50'd1771,50'd433},{50'd87,50'd508},{50'd1857,50'd1898},{50'd686,50'd84},{50'd1141,50'd1703},{50'd1394,50'd917},
        {50'd387,50'd1194},{50'd1594,50'd1183},{50'd724,50'd669},{50'd961,50'd1137},{50'd1171,50'd1045},{50'd1248,50'd1473},{50'd1975,50'd112},{50'd1075,50'd353},
        {50'd1676,50'd1576},{50'd1005,50'd1426},{50'd109,50'd1887},{50'd78,50'd455},{50'd1184,50'd2032},{50'd1256,50'd2024},{50'd770,50'd830},{50'd1044,50'd604},
        {50'd1790,50'd394},{50'd1591,50'd735},{50'd518,50'd261},{50'd201,50'd687},{50'd67,50'd1820},{50'd2013,50'd40},{50'd17,50'd195},{50'd1566,50'd1260},
        {50'd1569,50'd1843},{50'd1470,50'd1452},{50'd1989,50'd1233},{50'd1392,50'd1361},{50'd1696,50'd994},{50'd1847,50'd1110},{50'd1106,50'd537},{50'd668,50'd896},
        {50'd1229,50'd1366},{50'd1769,50'd263},{50'd137,50'd423},{50'd296,50'd1047},{50'd1715,50'd708},{50'd2030,50'd39},{50'd1891,50'd414},{50'd1855,50'd947},
        {50'd406,50'd1561},{50'd1352,50'd1035},{50'd565,50'd265},{50'd1996,50'd1701},{50'd91,50'd1236},{50'd1486,50'd395},{50'd583,50'd1580},{50'd95,50'd1711},
        {50'd1187,50'd1078},{50'd1360,50'd277},{50'd1446,50'd1648},{50'd1354,50'd1577},{50'd906,50'd461},{50'd664,50'd216},{50'd1132,50'd226},{50'd379,50'd1332},
        {50'd711,50'd1379},{50'd1928,50'd648},{50'd2016,50'd1865},{50'd1603,50'd637},{50'd816,50'd1315},{50'd1749,50'd480},{50'd24,50'd446},{50'd738,50'd1706},
        {50'd1814,50'd1791},{50'd466,50'd1050},{50'd1174,50'd158},{50'd160,50'd202},{50'd1060,50'd271},{50'd577,50'd791},{50'd1277,50'd1700},{50'd1010,50'd1323},
        {50'd1852,50'd1097},{50'd1270,50'd129},{50'd1529,50'd1056},{50'd992,50'd1027},{50'd59,50'd1513},{50'd674,50'd2022},{50'd933,50'd1369},{50'd576,50'd597},
        {50'd601,50'd644},{50'd1549,50'd852},{50'd697,50'd580},{50'd1871,50'd469},{50'd1375,50'd1949},{50'd1766,50'd1516},{50'd2004,50'd1310},{50'd598,50'd1937},
        {50'd234,50'd1794},{50'd1099,50'd76},{50'd372,50'd1383},{50'd99,50'd854},{50'd1890,50'd1761},{50'd855,50'd826},{50'd1609,50'd986},{50'd1826,50'd1475},
        {50'd925,50'd1640},{50'd894,50'd1325},{50'd1199,50'd915},{50'd38,50'd1147},{50'd1878,50'd203},{50'd2029,50'd730},{50'd1207,50'd1350},{50'd177,50'd1267},
        {50'd1424,50'd1707},{50'd1029,50'd219},{50'd1815,50'd424},{50'd188,50'd1746},{50'd506,50'd247},{50'd1262,50'd1977},{50'd996,50'd662},{50'd910,50'd661},
        {50'd793,50'd1610},{50'd589,50'd349},{50'd617,50'd113},{50'd36,50'd978},{50'd63,50'd180},{50'd243,50'd931},{50'd585,50'd1656},{50'd1764,50'd1850},
        {50'd882,50'd1157},{50'd1950,50'd1242},{50'd530,50'd1269},{50'd647,50'd504},{50'd456,50'd166},{50'd1278,50'd1122},{50'd1013,50'd559},{50'd1743,50'd542},
        {50'd2009,50'd827},{50'd1389,50'd1119},{50'd1586,50'd1875},{50'd374,50'd1434},{50'd1959,50'd1822},{50'd744,50'd972},{50'd1731,50'd689},{50'd1365,50'd775},
        {50'd1678,50'd13},{50'd893,50'd1213},{50'd1234,50'd1584},{50'd787,50'd795},{50'd1385,50'd1088},{50'd281,50'd800},{50'd1160,50'd863},{50'd352,50'd260},
        {50'd127,50'd774},{50'd1093,50'd1940},{50'd305,50'd2010},{50'd1291,50'd1779},{50'd413,50'd325},{50'd1778,50'd706},{50'd1240,50'd573},{50'd1844,50'd922},
        {50'd445,50'd1289},{50'd1927,50'd2028},{50'd536,50'd1338},{50'd399,50'd819},{50'd1564,50'd163},{50'd1614,50'd562},{50'd956,50'd1567},{50'd1422,50'd1956},
        {50'd982,50'd705},{50'd176,50'd510},{50'd289,50'd338},{50'd1806,50'd454},{50'd1899,50'd1300},{50'd1324,50'd1471},{50'd703,50'd1710},{50'd1118,50'd170},
        {50'd1105,50'd638},{50'd1643,50'd1512},{50'd320,50'd546},{50'd663,50'd1259},{50'd1388,50'd489},{50'd280,50'd1115},{50'd83,50'd96},{50'd1283,50'd1449},
        {50'd790,50'd1936},{50'd1997,50'd1873},{50'd1402,50'd574},{50'd810,50'd765},{50'd1727,50'd1028},{50'd732,50'd1395},{50'd867,50'd935},{50'd1428,50'd1382},
        {50'd673,50'd2025},{50'd1222,50'd435},{50'd1401,50'd511},{50'd1108,50'd1698},{50'd102,50'd1507},{50'd367,50'd1976},{50'd1983,50'd1930},{50'd1436,50'd1347},
        {50'd2045,50'd870},{50'd842,50'd135},{50'd983,50'd988},{50'd1348,50'd1808},{50'd1483,50'd1916},{50'd965,50'd579},{50'd1249,50'd1489},{50'd1602,50'd1635},
        {50'd1508,50'd588},{50'd1405,50'd1694},{50'd1776,50'd1720},{50'd501,50'd887},{50'd1203,50'd1345},{50'd1742,50'd756},{50'd1355,50'd1785},{50'd110,50'd238},
        {50'd1828,50'd1279},{50'd932,50'd1114},{50'd1903,50'd1672},{50'd1964,50'd400},{50'd1318,50'd1371},{50'd1178,50'd1535},{50'd1800,50'd1874},{50'd781,50'd297},
        {50'd1835,50'd2034},{50'd1819,50'd1931},{50'd1912,50'd1419},{50'd1195,50'd1902},{50'd868,50'd5},{50'd1824,50'd1113},{50'd1469,50'd377},{50'd250,50'd1510},
        {50'd295,50'd1070},{50'd331,50'd1440},{50'd1590,50'd1679},{50'd428,50'd1995},{50'd618,50'd1859},{50'd760,50'd1854},{50'd1180,50'd727},{50'd1686,50'd1443},
        {50'd1626,50'd118},{50'd1116,50'd1313},{50'd1214,50'd1667},{50'd979,50'd1172},{50'd482,50'd876},{50'd904,50'd1437},{50'd1782,50'd1464},{50'd709,50'd484},
        {50'd1476,50'd1265},{50'd1125,50'd1098},{50'd364,50'd797},{50'd616,50'd694},{50'd1144,50'd183},{50'd27,50'd1257},{50'd293,50'd1601},{50'd1420,50'd133},
        {50'd1339,50'd1103},{50'd1716,50'd582},{50'd523,50'd15},{50'd699,50'd1798},{50'd227,50'd52},{50'd1504,50'd2005},{50'd1723,50'd1525},{50'd1933,50'd1801},
        {50'd1043,50'd1637},{50'd35,50'd507},{50'd1169,50'd602},{50'd104,50'd1409},{50'd25,50'd245},{50'd794,50'd287},{50'd1168,50'd1768},{50'd1287,50'd1658},
        {50'd462,50'd1688},{50'd997,50'd1653},{50'd1210,50'd607},{50'd998,50'd1250},{50'd266,50'd1190},{50'd1458,50'd404},{50'd1986,50'd107},{50'd1729,50'd1336},
        {50'd595,50'd476},{50'd1605,50'd1528},{50'd1748,50'd1988},{50'd233,50'd208},{50'd993,50'd749},{50'd11,50'd73},{50'd859,50'd864},{50'd685,50'd1399},
        {50'd1935,50'd1496},{50'd926,50'd531},{50'd629,50'd493},{50'd1456,50'd108},{50'd1797,50'd393},{50'd1059,50'd298},{50'd1435,50'd952},{50'd779,50'd676},
        {50'd1812,50'd214},{50'd1929,50'd960},{50'd282,50'd1721},{50'd270,50'd452},{50'd1608,50'd716},{50'd1834,50'd554},{50'd513,50'd1223},{50'd1258,50'd1926},
        {50'd119,50'd268},{50'd1033,50'd339},{50'd164,50'd1284},{50'd801,50'd702},{50'd179,50'd903},{50'd1219,50'd715},{50'd957,50'd603},{50'd1718,50'd851},
        {50'd385,50'd1480},{50'd1290,50'd23},{50'd623,50'd1292},{50'd272,50'd0},{50'd1100,50'd909},{50'd1170,50'd953},{50'd1046,50'd999},{50'd683,50'd1671},
        {50'd1164,50'd653},{50'd628,50'd534},{50'd1616,50'd1090},{50'd103,50'd625},{50'd1900,50'd1705},{50'd1282,50'd1193},{50'd328,50'd1391},{50'd612,50'd757},
        {50'd1685,50'd1969},{50'd557,50'd1642},{50'd822,50'd1211},{50'd1307,50'd1582},{50'd1129,50'd970},{50'd390,50'd532},{50'd946,50'd141},{50'd4,50'd431},
        {50'd458,50'd165},{50'd813,50'd1955},{50'd1299,50'd1049},{50'd908,50'd1036},{50'd389,50'd581},{50'd1612,50'd1578},{50'd1534,50'd1911},{50'd985,50'd1531},
        {50'd1697,50'd981},{50'd1505,50'd1737},{50'd1281,50'd1433},{50'd359,50'd1726},{50'd1124,50'd145},{50'd1185,50'd199},{50'd1201,50'd2019},{50'd408,50'd420},
        {50'd1055,50'd360},{50'd564,50'd1632},{50'd1877,50'd1128},{50'd950,50'd1831},{50'd2003,50'd754},{50'd1682,50'd1560},{50'd371,50'd1934},{50'd1982,50'd1714},
        {50'd1666,50'd220},{50'd1619,50'd1359},{50'd350,50'd474},{50'd70,50'd1271},{50'd1818,50'd539},{50'd1625,50'd802},{50'd32,50'd1418},{50'd1408,50'd1495},
        {50'd1319,50'd449},{50'd86,50'd1568},{50'd290,50'd175},{50'd1488,50'd22},{50'd1331,50'd307},{50'd2027,50'd516},{50'd237,50'd278},{50'd789,50'd1398},
        {50'd1312,50'd1979},{50'd840,50'd1615},{50'd761,50'd1212},{50'd808,50'd670},{50'd373,50'd729},{50'd1427,50'd1139},{50'd1152,50'd1559},{50'd987,50'd680},
        {50'd596,50'd1487},{50'd1081,50'd1162},{50'd1762,50'd620},{50'd284,50'd1372},{50'd684,50'd1163},{50'd392,50'd873},{50'd1151,50'd69},{50'd88,50'd1973},
        {50'd440,50'd1880},{50'd899,50'd1096},{50'd1652,50'd1848},{50'd487,50'd2036},{50'd1004,50'd1544},{50'd386,50'd543},{50'd1455,50'd1337},{50'd417,50'd1941},
        {50'd1462,50'd190},{50'd1253,50'd122},{50'd1987,50'd1066},{50'd1386,50'd318},{50'd2041,50'd274},{50'd541,50'd593},{50'd447,50'd1981},{50'd905,50'd354},
        {50'd1241,50'd701},{50'd1370,50'd1574},{50'd1176,50'd1673},{50'd355,50'd1209},{50'd1773,50'd33},{50'd860,50'd1439},{50'd1189,50'd1235},{50'd1745,50'd898},
        {50'd1317,50'd1905},{50'd1509,50'd1647},{50'd878,50'd722},{50'd1681,50'd1868},{50'd1228,50'd1551},{50'd2002,50'd229},{50'd681,50'd928},{50'd384,50'd655},
        {50'd286,50'd1166},{50'd1491,50'd1406},{50'd486,50'd366},{50'd1984,50'd57},{50'd1073,50'd763},{50'd1669,50'd1811},{50'd1161,50'd1384},{50'd558,50'd1208},
        {50'd432,50'd1500},{50'd1003,50'd866},{50'd806,50'd892},{50'd1554,50'd448},{50'd427,50'd1344},{50'd1799,50'd914},{50'd470,50'd346},{50'd630,50'd1217},
        {50'd124,50'd679},{50'd1430,50'd1919},{50'd422,50'd75},{50'd526,50'd865},{50'd1943,50'd584},{50'd1205,50'd65},{50'd1895,50'd34},{50'd567,50'd1932},
        {50'd161,50'd1829},{50'd1126,50'd1804},{50'd1091,50'd248},{50'd54,50'd1639},{50'd938,50'd1553},{50'd242,50'd1650},{50'd1215,50'd441},{50'd1136,50'd627},
        {50'd936,50'd396},{50'd205,50'd1901},{50'd1111,50'd1008},{50'd174,50'd1583},{50'd734,50'd1477},{50'd1404,50'd1954},{50'd2047,50'd111},{50'd1074,50'd412},
        {50'd460,50'd1167},{50'd1546,50'd1381},{50'd1532,50'd919},{50'd1484,50'd321},{50'd306,50'd1368},{50'd1104,50'd1654},{50'd640,50'd51},{50'd236,50'd712},
        {50'd490,50'd570},{50'd189,50'd61},{50'd1474,50'd1674},{50'd1182,50'd1052},{50'd1668,50'd1837},{50'd478,50'd1465},{50'd147,50'd1225},{50'd138,50'd488},
        {50'd154,50'd1246},{50'd368,50'd1821},{50'd1751,50'd1951},{50'd693,50'd544},{50'd654,50'd1138},{50'd1813,50'd818},{50'd1565,50'd786},{50'd1273,50'd551},
        {50'd1305,50'd976},{50'd29,50'd740},{50'd241,50'd315},{50'd1879,50'd1396},{50'd173,50'd836},{50'd1467,50'd788},{50'd820,50'd943},{50'd1227,50'd592},
        {50'd881,50'd7},{50'd1341,50'd1712},{50'd416,50'd1897},{50'd741,50'd1866},{50'd1482,50'd857},{50'd512,50'd714},{50'd1886,50'd1695},{50'd1542,50'd94},
        {50'd1770,50'd1413},{50'd675,50'd1524},{50'd58,50'd2006},{50'd1841,50'd1094},{50'd401,50'd783},{50'd611,50'd1362},{50'd1380,50'd1025},{50'd101,50'd639},
        {50'd1085,50'd805},{50'd358,50'd323},{50'd1197,50'd1089},{50'd1781,50'd519},{50'd514,50'd1511},{50'd437,50'd733},{50'd157,50'd545},{50'd1340,50'd1054},
        {50'd1924,50'd1763},{50'd1758,50'd1888},{50'd1882,50'd77},{50'd930,50'd1077},{50'd1351,50'd1058},{50'd1947,50'd861},{50'd1102,50'd114},{50'd843,50'd1759},
        {50'd1518,50'd217},{50'd149,50'd249},{50'd890,50'd1015},{50'd1809,50'd1481},{50'd150,50'd182},{50'd1441,50'd768},{50'd657,50'd1757},{50'd148,50'd621},
        {50'd563,50'd1846},{50'd1067,50'd240},{50'd1244,50'd762},{50'd1072,50'd1177},{50'd1342,50'd505},{50'd1295,50'd1680},{50'd934,50'd376},{50'd746,50'd1552},
        {50'd615,50'd631},{50'd1689,50'd1883},{50'd1296,50'd6},{50'd751,50'd1889},{50'd184,50'd162},{50'd16,50'd1328},{50'd1068,50'd1453},{50'd1592,50'd1198},
        {50'd312,50'd1833},{50'd1699,50'd397},{50'd1810,50'd1173},{50'd1321,50'd844},{50'd944,50'd660},{50'd721,50'd209},{50'd1002,50'd50},{50'd60,50'd1744},
        {50'd308,50'd771},{50'd1991,50'd1308},{50'd856,50'd143},{50'd224,50'd954},{50'd1693,50'd921},{50'd707,50'd326},{50'd811,50'd1573},{50'd1142,50'd1376},
        {50'd8,50'd159},{50'd121,50'd1860},{50'd115,50'd2038},{50'd64,50'd1725},{50'd1537,50'd1514},{50'd257,50'd1521},{50'd1921,50'd1101},{50'd792,50'd831},
        {50'd1558,50'd838},{50'd1285,50'd600},{50'd425,50'd313},{50'd330,50'd1736},{50'd1020,50'd776},{50'd1061,50'd499},{50'd608,50'd535},{50'd324,50'd1238},
        {50'd1251,50'd1600},{50'd1550,50'd1123},{50'd1750,50'd1216},{50'd1179,50'd1738},{50'd28,50'd1175},{50'd1832,50'd465},{50'd2033,50'd1397},{50'd343,50'd969},
        {50'd1607,50'd450},{50'd1863,50'd1817},{50'd1472,50'd672},{50'd1675,50'd1760},{50'd571,50'd1254},{50'd1186,50'd759},{50'd1881,50'd941},{50'd273,50'd410},
        {50'd1031,50'd380},{50'd719,50'd995},{50'd2008,50'd951},{50'd1793,50'd1717},{50'd1356,50'd1970},{50'd677,50'd619},{50'd351,50'd847},{50'd464,50'd1918},
        {50'd1772,50'd743},{50'd303,50'd902},{50'd1021,50'd222},{50'd750,50'd144},{50'd90,50'd1306},{50'd971,50'd1353},{50'd1461,50'd1038},{50'd212,50'd329},
        {50'd889,50'd2031},{50'd1585,50'd1403},{50'd370,50'd1494},{50'd1611,50'd1303},{50'd1965,50'd503},{50'd927,50'd1084},{50'd736,50'd832},{50'd667,50'd1327},
        {50'd1107,50'd49},{50'd1322,50'd1499},{50'd2039,50'd920},{50'd1407,50'd197},{50'd89,50'd991},{50'd1631,50'd553},{50'd231,50'd649},{50'd1849,50'd635},
        {50'd1972,50'd1665},{50'd1011,50'd1649},{50'd973,50'd232},{50'd1133,50'd849},{50'd522,50'd1755},{50'd451,50'd43},{50'd1644,50'd1083},{50'd496,50'd1181},
        {50'd168,50'd720},{50'd335,50'd1786},{50'd1774,50'd210},{50'd1914,50'd463},{50'd1335,50'd1309},{50'd1006,50'd1827},{50'd1862,50'd1520},{50'd1906,50'd1007},
        {50'd524,50'd1953},{50'd605,50'd116},{50'd1836,50'd1358},{50'd1017,50'd1754},{50'd200,50'd610},{50'd875,50'd430},{50'd198,50'd883},{50'd136,50'd10},
        {50'd1624,50'd126},{50'd1709,50'd225},{50'd2011,50'd1204},{50'd1633,50'd1620},{50'd3,50'd1719},{50'd213,50'd1032},{50'd239,50'd2000},{50'd1266,50'd587},
        {50'd194,50'd1952},{50'd1272,50'd566},{50'd207,50'd812},{50'd737,50'd1670},{50'd769,50'd1206},{50'd2018,50'd178},{50'd1466,50'd169},{50'd186,50'd276},
        {50'd337,50'd578},{50'd1243,50'd509},{50'd1051,50'd1390},{50'd586,50'd723},{50'd1892,50'd1562},{50'd319,50'd1506},{50'd1343,50'd1053},{50'd911,50'd1450},
        {50'd1628,50'd1026},{50'd632,50'd45},{50'd989,50'd1885},{50'd798,50'd1651},{50'd652,50'd434},{50'd309,50'd1636},{50'd246,50'd1845},{50'd671,50'd106},
        {50'd645,50'd146},{50'd807,50'd529},{50'd1239,50'd409},{50'd1589,50'd1530},{50'd1459,50'd1226},{50'd1024,50'd1158},{50'd93,50'd1146},{50'd1065,50'd966},
        {50'd1076,50'd1445},{50'd1864,50'd411},{50'd1134,50'd1966},{50'd1998,50'd1030},{50'd80,50'd907},{50'd835,50'd877},{50'd1638,50'd185},{50'd1357,50'd1596},
        {50'd945,50'd294},{50'd888,50'd1330},{50'd171,50'd1942},{50'd1604,50'd1288},{50'd421,50'd569},{50'd1165,50'd1867},{50'd785,50'd624},{50'd1663,50'd363},
        {50'd1522,50'd1922},{50'd1816,50'd823},{50'd646,50'd803},{50'd1572,50'd916},{50'd302,50'd68},{50'd1830,50'd948},{50'd1961,50'd301},{50'd606,50'd1109},
        {50'd1159,50'd2},{50'd251,50'd923},{50'd1255,50'd1492},{50'd398,50'd267},{50'd18,50'd391},{50'd1264,50'd1618},{50'd895,50'd1872},{50'd1939,50'd1597},
        {50'd123,50'd1301},{50'd678,50'd967},{50'd495,50'd494},{50'd1948,50'd1747},{50'd1063,50'd651},{50'd1425,50'd407},{50'd1377,50'd357},{50'd42,50'd1784},
        {50'd884,50'd402},{50'd1765,50'd764},{50'd132,50'd340},{50'd650,50'd1415},{50'd1120,50'd26},{50'd1595,50'd1588},{50'd1218,50'd696},{50'd2020,50'd1634},
        {50'd1980,50'd1519},{50'd1730,50'd92},{50'd1498,50'd347},{50'd1451,50'd192},{50'd342,50'd814},{50'd1040,50'd959},{50'd853,50'd528},{50'd1095,50'd1796},
        {50'd140,50'd1735},{50'd869,50'd1329},{50'd1230,50'd1925},{50'd2026,50'd48},{50'd235,50'd262},{50'd1374,50'd172},{50'd1431,50'd327},{50'd2017,50'd1896},
        {50'd120,50'd1432},{50'd1022,50'd525},{50'd382,50'd142},{50'd1915,50'd47},{50'd2021,50'd1593},{50'd71,50'd1400},{50'd21,50'd1149},{50'd1231,50'd1807},
        {50'd1543,50'd291},{50'd1079,50'd990},{50'd1946,50'd825},{50'd1333,50'd1071},{50'd1460,50'd275},{50'd752,50'd1780},{50'd117,50'd1023},{50'd1293,50'd977},
        {50'd918,50'd1581},{50'd1838,50'd230},{50'd255,50'd1622},{50'd1188,50'd1662},{50'd1148,50'd1019},{50'd1014,50'd939},{50'd1547,50'd1092},{50'd218,50'd299},
        {50'd1704,50'd731},{50'd439,50'd1570},{50'd1967,50'd666},{50'd1908,50'd1286},{50'd1468,50'd1690},{50'd1393,50'd549},{50'd984,50'd1001},{50'd453,50'd1555},
        {50'd1753,50'd1224},{50'd256,50'd2014},{50'd1938,50'd356},{50'd471,50'd1920},{50'd369,50'd472},{50'd1200,50'd1621},{50'd1739,50'd758},{50'd1788,50'd862},
        {50'd1153,50'd891},{50'd913,50'd572},{50'd1805,50'd1733},{50'd912,50'd590},{50'd477,50'd1298},{50'd897,50'd457},{50'd656,50'd300},{50'd500,50'd139},
        {50'd974,50'd2042},{50'd443,50'd9},{50'd436,50'd829},{50'd766,50'd634},{50'd1575,50'd1485},{50'd1907,50'd796},{50'd1740,50'd874},{50'd85,50'd167},
        {50'd1117,50'd426},{50'd691,50'd31},{50'd533,50'd2023},{50'd886,50'd283},{50'd599,50'd690},{50'd481,50'd1909},{50'd1692,50'd880},{50'd497,50'd1993},
        {50'd622,50'd772},{50'd748,50'd1630},{50'd1221,50'd1448},{50'd665,50'd403},{50'd1062,50'd1131},{50'd521,50'd942},{50'd1839,50'd1557},{50'd1302,50'd1490},
        {50'd1478,50'd19},{50'd1143,50'd556},{50'd1039,50'd964},{50'd181,50'd552},{50'd1533,50'd334},{50'd828,50'd739},{50'd1527,50'd74},{50'd1252,50'd1861},
        {50'd1,50'd2046},{50'd1853,50'd362},{50'd1412,50'd1958},{50'd473,50'd1884},{50'd626,50'd1416},{50'd1893,50'd485},{50'd975,50'd1598},{50'd1274,50'd1304},
        {50'd594,50'd1130},{50'd924,50'd310},{50'd20,50'd1994},{50'd1156,50'd717},{50'd2012,50'd1276},{50'd742,50'd782},{50'd130,50'd777},{50'd614,50'd688},
        {50'd438,50'd1438},{50'd540,50'd79},{50'd799,50'd1775},{50'd1429,50'd833},{50'd254,50'd745},{50'd560,50'd1606},{50'd704,50'd1155},{50'd152,50'd1501},
        {50'd98,50'd378},{50'd1275,50'd1587},{50'd1263,50'd1540},{50'd1363,50'd1985},{50'd317,50'd1541},{50'd336,50'd1414},{50'd710,50'd1823},{50'd718,50'd1978},
        {50'd1783,50'd259},{50'd316,50'd1563},{50'd475,50'd846},{50'd1373,50'd228},{50'd613,50'd269},{50'd1346,50'd1064},{50'd1121,50'd1913},{50'd520,50'd223},
        {50'd12,50'd37},{50'd1387,50'd467},{50'd1314,50'd66},{50'd322,50'd1856},{50'd53,50'd134},{50'd809,50'd1000},{50'd968,50'd187},{50'd1140,50'd1945},
        {50'd848,50'd1545},{50'd1870,50'd1645},{50'd1992,50'd1974},{50'd1722,50'd1802},{50'd1247,50'd279},{50'd824,50'd834},{50'd1220,50'd1687},{50'd418,50'd698},
        {50'd1752,50'd1655},{50'd900,50'd444},{50'd1261,50'd2043},{50'd962,50'd1660},{50'd728,50'd285},{50'd1421,50'd1497},{50'd1990,50'd1999},{50'd1617,50'd1297},
        {50'd1069,50'd858},{50'd193,50'd845},{50'd817,50'd1792},{50'd515,50'd1526},{50'd568,50'd1517},{50'd1613,50'd2015},{50'd498,50'd1150},{50'd191,50'd538},
        {50'd2007,50'd206},{50'd1191,50'd1691},{50'd1457,50'd1311},{50'd850,50'd1728},{50'd1237,50'd1963},{50'd1661,50'd125},{50'd468,50'd30},{50'd1756,50'd1657},
        {50'd1145,50'd1627},{50'd633,50'd1057},{50'd383,50'd365},{50'd1320,50'd215},{50'd747,50'd483},{50'd937,50'd1910},{50'd1479,50'd949},{50'd502,50'd131},
        {50'd2037,50'd55},{50'd1154,50'd1548},{50'd1280,50'd2001},{50'd211,50'd841},{50'd1042,50'd1493},{50'd1080,50'd62},{50'd492,50'd304},{50'd1917,50'd821},
        {50'd753,50'd1579},{50'd1202,50'd1536},{50'd682,50'd1539},{50'd82,50'd804},{50'd1732,50'd81},{50'd1444,50'd879},{50'd1112,50'd1018},{50'd288,50'd361},
        {50'd344,50'd1842},{50'd388,50'd1048},{50'd1659,50'd778},{50'd755,50'd1777},{50'd97,50'd901},{50'd726,50'd837},{50'd1571,50'd1683},{50'd253,50'd871},
        {50'd1127,50'd1708},{50'd1641,50'd658},{50'd1232,50'd258},{50'd591,50'd1734},{50'd955,50'd1858},{50'd1523,50'd156},{50'd1869,50'd1795},{50'd659,50'd1463},
        {50'd1411,50'd1556},{50'd1538,50'd1724},{50'd1245,50'd527},{50'd292,50'd244},{50'd1876,50'd153},{50'd1971,50'd415},{50'd767,50'd1378},{50'd963,50'd1787},
        {50'd1825,50'd491},{50'd885,50'd547},{50'd1629,50'd1664},{50'd442,50'd2035},{50'd1268,50'd784},{50'd773,50'd1423},{50'd196,50'd1960},{50'd41,50'd44}};



end


//read
always @ ( posedge clk )
begin
    if (en)
        dob <= ram[addrb];
end


//write
always @ (posedge clk)
begin
    if (we && en)
        ram[addra] <= dia;
end

endmodule
